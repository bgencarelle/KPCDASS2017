// adc_test.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module adc_test (
		input  wire        adc_pll_clock_clk,          //    adc_pll_clock.clk
		input  wire        adc_pll_locked_export,      //   adc_pll_locked.export
		input  wire        clock_clk,                  //            clock.clk
		input  wire        reset_sink_reset_n,         //       reset_sink.reset_n
		input  wire [6:0]  sample_store_csr_address,   // sample_store_csr.address
		input  wire        sample_store_csr_read,      //                 .read
		input  wire        sample_store_csr_write,     //                 .write
		input  wire [31:0] sample_store_csr_writedata, //                 .writedata
		output wire [31:0] sample_store_csr_readdata,  //                 .readdata
		output wire        sample_store_irq_irq,       // sample_store_irq.irq
		input  wire        sequencer_csr_address,      //    sequencer_csr.address
		input  wire        sequencer_csr_read,         //                 .read
		input  wire        sequencer_csr_write,        //                 .write
		input  wire [31:0] sequencer_csr_writedata,    //                 .writedata
		output wire [31:0] sequencer_csr_readdata      //                 .readdata
	);

	adc_test_modular_dual_adc_0 modular_dual_adc_0 (
		.clock_clk                  (clock_clk),                  //            clock.clk
		.reset_sink_reset_n         (reset_sink_reset_n),         //       reset_sink.reset_n
		.adc_pll_clock_clk          (adc_pll_clock_clk),          //    adc_pll_clock.clk
		.adc_pll_locked_export      (adc_pll_locked_export),      //   adc_pll_locked.export
		.sequencer_csr_address      (sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       (sample_store_irq_irq)        // sample_store_irq.irq
	);

endmodule
