
module issp (
	source);	

	output	[0:0]	source;
endmodule
