module midi_input (
input wire note_on,
input wire [6:0] note_number,
input wire note_off,
input wire velocity,
input wire pitch
);

endmodule