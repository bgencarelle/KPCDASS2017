
module clock_buff (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
